-- CPU
library IEEE;
library WORK;

use IEEE.STD_LOGIC_1164.all;
use IEEE.numeric_std.all;
use WORK.CPU_LIB.all;

entity CPU is
  port
    (
    -- Input ports
      clk		: STD_LOGIC;
--    reset		: STD_LOGIC;
--    load 		: STD_LOGIC;
--    stall 	: STD_LOGIC;

		-- Output ports	
    );
end CPU;

architecture arch of CPU is

begin	
end arch;